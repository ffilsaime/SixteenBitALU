/* ALU unit gate delay simulation used ot determine the average delay
*/

/* ALU unit gate delay simulation used to determine temporal delays
*/

/*
ALU zero delay simulation
*/

// this is the full adder for alu
`timescale 1ns/1ns
module fulladder(a,b,c,s,cout);
input a,b,c;
output s, cout;
wire axorb, bandc, canda, aandb; 
xor #1
    z1(axorb, a, b),
    z2(s, axorb, c);
and #1
    z3(bandc, b, c),
    z4(canda, c, a),
    z5(aandb, a, b);
or #1
    z6(cout, bandc, canda, aandb);
endmodule 

//2 to 1 mux
`timescale 1ns/1ns
module twotoone(first, second, select, choice);
input first, second, select;
output choice;
wire fsel, ssel, notsel;

not #1 y1(notsel, select);
and #1 y2(fsel, first, notsel);
and #1 y3(ssel, second, select);
or #1 y4(choice, ssel, fsel);
endmodule

//4 to 1 mux
`timescale 1ns/1ns
module fourToOne(sel, sel2, zero, one, two, three, selected);
input sel, sel2, zero, one, two, three;
output selected;
wire notsel, notsel2, w1, w2, w3, w4;

not #1
    x0(notsel, sel),
    x1(notsel2, sel2);
and #1 x2(w1, zero, notsel2, notsel);
and #1 x3(w2, two, sel, notsel2);
and #1 x4(w3, one, notsel, sel2);
and #1 x5(w4, three, sel2, sel);
or #1 x6(selected, w1, w2, w3, w4);
endmodule

//this is a 1 bit alu 
`timescale 1ns/1ns
module onealu(a, b, cin, s, cout, less, op, choice,q);
input a, b, cin, less; 
input [2:0] op;
output s, cout, choice, q;
wire aandb, aorb, notb;

not #1 t6(notb, b);
and #1 t5(aandb,a,b); // the and operation
or #1 t4(aorb, a,b); // the or operation
twotoone t1(b, notb, op[2], choice); // creates the 2 to 1 mux
fulladder t2(a, choice, cin, s, cout); // the adder of the alu
fourToOne t3(op[1], op[0], aandb, aorb, s, less, q);
endmodule

// this is the full alu
module sixteenBitalu(a, b, s, cout, op, choice, q);
input [15:0] a, b;
input [2:0] op;
output [15:0] s, choice, c, q;
output cout;

onealu o1(a[0], b[0], op[2], s[0], c[0], s[15], op, choice[0],q[0]);
onealu o2(a[1], b[1], c[0], s[1], c[1], 0, op, choice[1],q[1]);
onealu o3(a[2], b[2], c[1], s[2], c[2], 0, op, choice[2], q[2]);
onealu o4(a[3], b[3], c[2], s[3], c[3], 0, op, choice[3], q[3]);

onealu o5(a[4], b[4], c[3], s[4], c[4], 0, op, choice[4], q[4]);
onealu o6(a[5], b[5], c[4], s[5], c[5], 0, op, choice[5], q[5]);
onealu o7(a[6], b[6], c[5], s[6], c[6], 0, op, choice[6], q[6]);
onealu o8(a[7], b[7], c[6], s[7], c[7], 0, op, choice[7], q[7]);

onealu o9(a[8], b[8], c[7], s[8], c[8], 0, op, choice[8], q[8]);
onealu o10(a[9], b[9], c[8], s[9], c[9], 0, op, choice[9], q[9]);
onealu o11(a[10], b[10], c[9], s[10], c[10], 0, op, choice[10], q[10]);
onealu o12(a[11], b[11], c[10], s[11], c[11], 0, op, choice[11], q[11]);

onealu o13(a[12], b[12], c[11], s[12], c[12], 0, op, choice[12], q[12]);
onealu o14(a[13], b[13], c[12], s[13], c[13], 0, op, choice[13], q[13]);
onealu o15(a[14], b[14], c[13], s[14], c[14], 0, op, choice[14], q[14]);
onealu o16(a[15], b[15], c[14], s[15], cout, 0, op, choice[15], q[15]);
endmodule

//the grand testbench for the 1000 inputs
`timescale 1ns/1ns
module testbench();
output reg [15:0] a, b;
output reg [2:0] op;
input [15:0] s, choice, q;
input cout;
sixteenBitalu s1(a, b, s, cout, op, choice, q);
initial
  begin
  $monitor($time,, "a=%d, b=%d, s=%d, cout=%b, op=%b, choice=%b, q=%d", a, b, s, cout, op, choice, q);
  $display($time,, "a=%d, b=%d, s=%d, cout=%b, op=%b, choice=%b, q=%d", a, b, s, cout, op, choice, q);
#30 a = 37215; b = 41581; op = 110;
#30 a = 50452; b = 40665; op = 110;
#30 a = 16435; b = 36713; op = 110;
#30 a = 1362; b = 29513; op = 110;
#30 a = 59893; b = 13238; op = 110;
#30 a = 38907; b = 44144; op = 110;
#30 a = 28931; b = 20459; op = 110;
#30 a = 53455; b = 43036; op = 110;
#30 a = 34099; b = 20682; op = 110;
#30 a = 49218; b = 38146; op = 110;
#30 a = 14738; b = 42682; op = 110;
#30 a = 59115; b = 26883; op = 110;
#30 a = 4457; b = 18500; op = 110;
#30 a = 54876; b = 28186; op = 110;
#30 a = 4156; b = 41607; op = 110;
#30 a = 45420; b = 36484; op = 110;
#30 a = 15725; b = 10904; op = 110;
#30 a = 48879; b = 33932; op = 110;
#30 a = 16221; b = 35641; op = 110;
#30 a = 34503; b = 22707; op = 110;
#30 a = 46259; b = 49780; op = 110;
#30 a = 32852; b = 26489; op = 110;
#30 a = 7893; b = 19413; op = 110;
#30 a = 58663; b = 22570; op = 110;
#30 a = 48210; b = 57602; op = 110;
#30 a = 31060; b = 47208; op = 110;
#30 a = 19330; b = 49783; op = 110;
#30 a = 28198; b = 42224; op = 110;
#30 a = 43301; b = 21282; op = 110;
#30 a = 11948; b = 31532; op = 110;
#30 a = 43368; b = 53464; op = 110;
#30 a = 35249; b = 35477; op = 110;
#30 a = 11719; b = 36210; op = 110;
#30 a = 37289; b = 43042; op = 110;
#30 a = 17484; b = 19303; op = 110;
#30 a = 20967; b = 46193; op = 110;
#30 a = 47285; b = 44519; op = 110;
#30 a = 29964; b = 29329; op = 110;
#30 a = 41204; b = 14610; op = 110;
#30 a = 42779; b = 57738; op = 110;
#30 a = 7696; b = 48435; op = 110;
#30 a = 15367; b = 56297; op = 110;
#30 a = 37320; b = 51004; op = 110;
#30 a = 34893; b = 55148; op = 110;
#30 a = 7064; b = 18271; op = 110;
#30 a = 13310; b = 52262; op = 110;
#30 a = 52180; b = 13254; op = 110;
#30 a = 4021; b = 1872; op = 110;
#30 a = 13457; b = 7119; op = 110;
#30 a = 23783; b = 7149; op = 110;
#30 a = 3267; b = 45096; op = 110;
#30 a = 36728; b = 31672; op = 110;
#30 a = 32353; b = 59331; op = 110;
#30 a = 48393; b = 40843; op = 110;
#30 a = 37253; b = 11958; op = 110;
#30 a = 9967; b = 33454; op = 110;
#30 a = 7535; b = 58834; op = 110;
#30 a = 33152; b = 51611; op = 110;
#30 a = 15561; b = 8925; op = 110;
#30 a = 21863; b = 17930; op = 110;
#30 a = 27749; b = 27310; op = 110;
#30 a = 41623; b = 31550; op = 110;
#30 a = 59395; b = 57604; op = 110;
#30 a = 28475; b = 30155; op = 110;
#30 a = 55311; b = 45796; op = 110;
#30 a = 45772; b = 13954; op = 110;
#30 a = 39591; b = 36014; op = 110;
#30 a = 41244; b = 5818; op = 110;
#30 a = 23674; b = 42747; op = 110;
#30 a = 51727; b = 16541; op = 110;
#30 a = 17771; b = 56596; op = 110;
#30 a = 37225; b = 38796; op = 110;
#30 a = 22421; b = 23410; op = 110;
#30 a = 1122; b = 37040; op = 110;
#30 a = 30088; b = 44141; op = 110;
#30 a = 2454; b = 24446; op = 110;
#30 a = 3538; b = 42659; op = 110;
#30 a = 17946; b = 30310; op = 110;
#30 a = 8506; b = 42984; op = 110;
#30 a = 34985; b = 43000; op = 110;
#30 a = 8677; b = 29540; op = 110;
#30 a = 10364; b = 33748; op = 110;
#30 a = 2459; b = 53838; op = 110;
#30 a = 54680; b = 38605; op = 110;
#30 a = 22755; b = 54499; op = 110;
#30 a = 22208; b = 43992; op = 110;
#30 a = 38411; b = 12130; op = 110;
#30 a = 21611; b = 18135; op = 110;
#30 a = 17476; b = 43783; op = 110;
#30 a = 34897; b = 44636; op = 110;
#30 a = 3754; b = 48386; op = 110;
#30 a = 30464; b = 33692; op = 110;
#30 a = 9890; b = 12819; op = 110;
#30 a = 23627; b = 38675; op = 110;
#30 a = 13724; b = 15141; op = 110;
#30 a = 28129; b = 55245; op = 110;
#30 a = 55255; b = 25348; op = 110;
#30 a = 35739; b = 57912; op = 110;
#30 a = 54147; b = 11228; op = 110;
#30 a = 43087; b = 44708; op = 110;
#30 a = 19970; b = 10255; op = 110;
#30 a = 12290; b = 56339; op = 110;
#30 a = 52168; b = 21331; op = 110;
#30 a = 52795; b = 3331; op = 110;
#30 a = 50370; b = 582; op = 110;
#30 a = 30482; b = 54773; op = 110;
#30 a = 5555; b = 16398; op = 110;
#30 a = 21607; b = 51769; op = 110;
#30 a = 23033; b = 5682; op = 110;
#30 a = 6158; b = 58232; op = 110;
#30 a = 47885; b = 3758; op = 110;
#30 a = 17128; b = 59005; op = 110;
#30 a = 42505; b = 1783; op = 110;
#30 a = 33710; b = 49089; op = 110;
#30 a = 48453; b = 37004; op = 110;
#30 a = 47846; b = 32531; op = 110;
#30 a = 9050; b = 28116; op = 110;
#30 a = 9176; b = 29344; op = 110;
#30 a = 29927; b = 13658; op = 110;
#30 a = 7066; b = 23652; op = 110;
#30 a = 28274; b = 13410; op = 110;
#30 a = 14184; b = 15373; op = 110;
#30 a = 17254; b = 1895; op = 110;
#30 a = 4623; b = 32391; op = 110;
#30 a = 13754; b = 24722; op = 110;
#30 a = 52328; b = 42122; op = 110;
#30 a = 29459; b = 32953; op = 110;
#30 a = 38434; b = 35549; op = 110;
#30 a = 54048; b = 20114; op = 110;
#30 a = 42456; b = 57573; op = 110;
#30 a = 39554; b = 11026; op = 110;
#30 a = 46722; b = 18894; op = 110;
#30 a = 53999; b = 6246; op = 110;
#30 a = 30407; b = 32884; op = 110;
#30 a = 38316; b = 58029; op = 110;
#30 a = 55727; b = 18638; op = 110;
#30 a = 52695; b = 45712; op = 110;
#30 a = 9975; b = 20024; op = 110;
#30 a = 3591; b = 46879; op = 110;
#30 a = 22206; b = 30460; op = 110;
#30 a = 49931; b = 48874; op = 110;
#30 a = 12636; b = 27773; op = 110;
#30 a = 44815; b = 20632; op = 110;
#30 a = 8883; b = 44671; op = 110;
#30 a = 606; b = 40871; op = 110;
#30 a = 33021; b = 5718; op = 110;
#30 a = 5377; b = 10625; op = 110;
#30 a = 24581; b = 29577; op = 110;
#30 a = 55269; b = 27800; op = 110;
#30 a = 43377; b = 24098; op = 110;
#30 a = 42106; b = 29566; op = 110;
#30 a = 22237; b = 44918; op = 110;
#30 a = 11863; b = 5027; op = 110;
#30 a = 51651; b = 35980; op = 110;
#30 a = 37083; b = 22347; op = 110;
#30 a = 16150; b = 17675; op = 110;
#30 a = 2063; b = 48843; op = 110;
#30 a = 13135; b = 45988; op = 110;
#30 a = 17032; b = 22880; op = 110;
#30 a = 31486; b = 33529; op = 110;
#30 a = 58472; b = 18733; op = 110;
#30 a = 15298; b = 45864; op = 110;
#30 a = 23747; b = 13807; op = 110;
#30 a = 26675; b = 27417; op = 110;
#30 a = 10239; b = 49566; op = 110;
#30 a = 21308; b = 38496; op = 110;
#30 a = 29205; b = 14306; op = 110;
#30 a = 2791; b = 24334; op = 110;
#30 a = 28149; b = 15183; op = 110;
#30 a = 1489; b = 5626; op = 110;
#30 a = 22630; b = 31391; op = 110;
#30 a = 58684; b = 44040; op = 110;
#30 a = 48490; b = 43595; op = 110;
#30 a = 49219; b = 27828; op = 110;
#30 a = 37247; b = 23430; op = 110;
#30 a = 31656; b = 8509; op = 110;
#30 a = 30402; b = 40245; op = 110;
#30 a = 55753; b = 9937; op = 110;
#30 a = 26575; b = 8591; op = 110;
#30 a = 12530; b = 720; op = 110;
#30 a = 42147; b = 56141; op = 110;
#30 a = 4908; b = 8383; op = 110;
#30 a = 25730; b = 35309; op = 110;
#30 a = 2962; b = 29548; op = 110;
#30 a = 51413; b = 14953; op = 110;
#30 a = 55460; b = 37849; op = 110;
#30 a = 36843; b = 49231; op = 110;
#30 a = 51668; b = 3175; op = 110;
#30 a = 14560; b = 16797; op = 110;
#30 a = 41566; b = 47969; op = 110;
#30 a = 15131; b = 55452; op = 110;
#30 a = 24309; b = 37377; op = 110;
#30 a = 44977; b = 20694; op = 110;
#30 a = 40184; b = 45250; op = 110;
#30 a = 19527; b = 42772; op = 110;
#30 a = 32260; b = 50180; op = 110;
#30 a = 15892; b = 36056; op = 110;
#30 a = 31555; b = 31830; op = 110;
#30 a = 35557; b = 42003; op = 110;
#30 a = 8706; b = 27299; op = 110;
#30 a = 14427; b = 23109; op = 110;
#30 a = 6016; b = 25563; op = 110;
#30 a = 3535; b = 10927; op = 110;
#30 a = 13730; b = 18109; op = 110;
#30 a = 56757; b = 53430; op = 110;
#30 a = 44835; b = 36798; op = 110;
#30 a = 10270; b = 57623; op = 110;
#30 a = 58697; b = 12696; op = 110;
#30 a = 1911; b = 21921; op = 110;
#30 a = 31859; b = 16594; op = 110;
#30 a = 7151; b = 23347; op = 110;
#30 a = 30926; b = 12456; op = 110;
#30 a = 534; b = 16147; op = 110;
#30 a = 999; b = 28951; op = 110;
#30 a = 42529; b = 10120; op = 110;
#30 a = 35195; b = 37383; op = 110;
#30 a = 39882; b = 50069; op = 110;
#30 a = 11305; b = 47733; op = 110;
#30 a = 58389; b = 43443; op = 110;
#30 a = 24457; b = 23580; op = 110;
#30 a = 19149; b = 20137; op = 110;
#30 a = 5815; b = 36160; op = 110;
#30 a = 42540; b = 27915; op = 110;
#30 a = 15879; b = 14582; op = 110;
#30 a = 15961; b = 16716; op = 110;
#30 a = 40092; b = 1683; op = 110;
#30 a = 50668; b = 38369; op = 110;
#30 a = 13428; b = 54960; op = 110;
#30 a = 40557; b = 5043; op = 110;
#30 a = 10331; b = 1559; op = 110;
#30 a = 53627; b = 52160; op = 110;
#30 a = 20960; b = 25644; op = 110;
#30 a = 47592; b = 33935; op = 110;
#30 a = 38308; b = 42971; op = 110;
#30 a = 6273; b = 5391; op = 110;
#30 a = 3694; b = 19642; op = 110;
#30 a = 27500; b = 58315; op = 110;
#30 a = 56220; b = 16666; op = 110;
#30 a = 54346; b = 9771; op = 110;
#30 a = 18517; b = 2032; op = 110;
#30 a = 15836; b = 1322; op = 110;
#30 a = 57049; b = 29370; op = 110;
#30 a = 9313; b = 24688; op = 110;
#30 a = 6489; b = 25552; op = 110;
#30 a = 31933; b = 15020; op = 110;
#30 a = 47363; b = 30953; op = 110;
#30 a = 37494; b = 41967; op = 110;
#30 a = 48918; b = 21735; op = 110;
#30 a = 16792; b = 19591; op = 110;
#30 a = 16180; b = 3968; op = 110;
#30 a = 11257; b = 1942; op = 110;
#30 a = 8021; b = 31082; op = 110;
#30 a = 10166; b = 8239; op = 110;
#30 a = 34808; b = 418; op = 110;
#30 a = 59131; b = 1549; op = 110;
#30 a = 22357; b = 54520; op = 110;
#30 a = 45218; b = 34512; op = 110;
#30 a = 2958; b = 12987; op = 110;
#30 a = 32723; b = 43541; op = 110;
#30 a = 43075; b = 38845; op = 110;
#30 a = 12362; b = 52976; op = 110;
#30 a = 31524; b = 13666; op = 110;
#30 a = 12983; b = 37257; op = 110;
#30 a = 3649; b = 18186; op = 110;
#30 a = 14302; b = 24080; op = 110;
#30 a = 48798; b = 41753; op = 110;
#30 a = 53854; b = 12958; op = 110;
#30 a = 5858; b = 36128; op = 110;
#30 a = 23951; b = 27817; op = 110;
#30 a = 9679; b = 32585; op = 110;
#30 a = 47172; b = 45636; op = 110;
#30 a = 54636; b = 42052; op = 110;
#30 a = 37169; b = 46673; op = 110;
#30 a = 41565; b = 30089; op = 110;
#30 a = 22150; b = 4036; op = 110;
#30 a = 29300; b = 21065; op = 110;
#30 a = 36441; b = 13301; op = 110;
#30 a = 33025; b = 37110; op = 110;
#30 a = 56705; b = 39777; op = 110;
#30 a = 22853; b = 21547; op = 110;
#30 a = 17662; b = 6686; op = 110;
#30 a = 50340; b = 36185; op = 110;
#30 a = 42871; b = 7097; op = 110;
#30 a = 37049; b = 55568; op = 110;
#30 a = 21339; b = 35086; op = 110;
#30 a = 53539; b = 40166; op = 110;
#30 a = 39529; b = 40707; op = 110;
#30 a = 32285; b = 43847; op = 110;
#30 a = 41451; b = 57218; op = 110;
#30 a = 2124; b = 53689; op = 110;
#30 a = 31901; b = 59761; op = 110;
#30 a = 28369; b = 58826; op = 110;
#30 a = 48524; b = 29039; op = 110;
#30 a = 10494; b = 22360; op = 110;
#30 a = 27897; b = 24365; op = 110;
#30 a = 52229; b = 53885; op = 110;
#30 a = 9532; b = 36358; op = 110;
#30 a = 16428; b = 18166; op = 110;
#30 a = 41637; b = 40221; op = 110;
#30 a = 40253; b = 16686; op = 110;
#30 a = 28094; b = 34386; op = 110;
#30 a = 24570; b = 52427; op = 110;
#30 a = 10093; b = 53792; op = 110;
#30 a = 43534; b = 20757; op = 110;
#30 a = 36054; b = 52950; op = 110;
#30 a = 47966; b = 29886; op = 110;
#30 a = 46908; b = 56943; op = 110;
#30 a = 21470; b = 31859; op = 110;
#30 a = 46056; b = 4945; op = 110;
#30 a = 47008; b = 21309; op = 110;
#30 a = 39586; b = 23871; op = 110;
#30 a = 45607; b = 6356; op = 110;
#30 a = 19900; b = 25595; op = 110;
#30 a = 31001; b = 10657; op = 110;
#30 a = 19791; b = 17756; op = 110;
#30 a = 33747; b = 33838; op = 110;
#30 a = 25885; b = 22631; op = 110;
#30 a = 16599; b = 46637; op = 110;
#30 a = 24981; b = 55469; op = 110;
#30 a = 10945; b = 5506; op = 110;
#30 a = 4596; b = 49217; op = 110;
#30 a = 44311; b = 5229; op = 110;
#30 a = 9449; b = 59508; op = 110;
#30 a = 11230; b = 24248; op = 110;
#30 a = 26001; b = 54255; op = 110;
#30 a = 38921; b = 19193; op = 110;
#30 a = 14241; b = 19212; op = 110;
#30 a = 53773; b = 43140; op = 110;
#30 a = 30498; b = 10738; op = 110;
#30 a = 32400; b = 45201; op = 110;
#30 a = 43095; b = 25131; op = 110;
#30 a = 18751; b = 3973; op = 110;
#30 a = 27162; b = 8451; op = 110;
#30 a = 31359; b = 11840; op = 110;
#30 a = 35428; b = 3807; op = 110;
#30 a = 39867; b = 13954; op = 110;
#30 a = 37675; b = 12152; op = 110;
#30 a = 16316; b = 27642; op = 110;
#30 a = 5893; b = 14611; op = 110;
#30 a = 11191; b = 21389; op = 110;
#30 a = 54443; b = 55582; op = 110;
#30 a = 46879; b = 33247; op = 110;
#30 a = 18553; b = 8; op = 110;
#30 a = 31388; b = 15682; op = 110;
#30 a = 25010; b = 56958; op = 110;
#30 a = 11540; b = 20888; op = 110;
#30 a = 59745; b = 34878; op = 110;
#30 a = 12389; b = 15142; op = 110;
#30 a = 3994; b = 47642; op = 110;
#30 a = 25332; b = 8855; op = 110;
#30 a = 57086; b = 17098; op = 110;
#30 a = 42784; b = 21353; op = 110;
#30 a = 22110; b = 49102; op = 110;
#30 a = 48240; b = 58969; op = 110;
#30 a = 26006; b = 36959; op = 110;
#30 a = 54187; b = 34630; op = 110;
#30 a = 44827; b = 7985; op = 110;
#30 a = 50566; b = 40388; op = 110;
#30 a = 19055; b = 26568; op = 110;
#30 a = 12599; b = 18112; op = 110;
#30 a = 39857; b = 26003; op = 110;
#30 a = 27529; b = 42347; op = 110;
#30 a = 42834; b = 39913; op = 110;
#30 a = 41416; b = 26181; op = 110;
#30 a = 40225; b = 38910; op = 110;
#30 a = 51516; b = 4679; op = 110;
#30 a = 1065; b = 22498; op = 110;
#30 a = 39891; b = 52460; op = 110;
#30 a = 4944; b = 7319; op = 110;
#30 a = 1911; b = 8381; op = 110;
#30 a = 47808; b = 910; op = 110;
#30 a = 48639; b = 42456; op = 110;
#30 a = 21123; b = 8061; op = 110;
#30 a = 47264; b = 6556; op = 110;
#30 a = 47687; b = 27998; op = 110;
#30 a = 53796; b = 58516; op = 110;
#30 a = 13473; b = 26758; op = 110;
#30 a = 22547; b = 34781; op = 110;
#30 a = 18349; b = 52672; op = 110;
#30 a = 174; b = 54102; op = 110;
#30 a = 39348; b = 30406; op = 110;
#30 a = 41307; b = 26755; op = 110;
#30 a = 58662; b = 33467; op = 110;
#30 a = 17593; b = 2046; op = 110;
#30 a = 50759; b = 44616; op = 110;
#30 a = 59829; b = 55515; op = 110;
#30 a = 40518; b = 16754; op = 110;
#30 a = 29974; b = 46645; op = 110;
#30 a = 5992; b = 28852; op = 110;
#30 a = 39827; b = 35898; op = 110;
#30 a = 11972; b = 47071; op = 110;
#30 a = 5061; b = 9489; op = 110;
#30 a = 23335; b = 5034; op = 110;
#30 a = 16055; b = 3555; op = 110;
#30 a = 34999; b = 4887; op = 110;
#30 a = 121; b = 7117; op = 110;
#30 a = 30165; b = 48291; op = 110;
#30 a = 24691; b = 18944; op = 110;
#30 a = 55964; b = 12169; op = 110;
#30 a = 1207; b = 49267; op = 110;
#30 a = 24806; b = 10037; op = 110;
#30 a = 2287; b = 1766; op = 110;
#30 a = 56589; b = 33024; op = 110;
#30 a = 40086; b = 50515; op = 110;
#30 a = 19406; b = 31597; op = 110;
#30 a = 35618; b = 57971; op = 110;
#30 a = 2314; b = 17566; op = 110;
#30 a = 19711; b = 29131; op = 110;
#30 a = 30663; b = 17940; op = 110;
#30 a = 38263; b = 41649; op = 110;
#30 a = 2964; b = 38753; op = 110;
#30 a = 18189; b = 38078; op = 110;
#30 a = 22889; b = 48939; op = 110;
#30 a = 19882; b = 57234; op = 110;
#30 a = 11180; b = 20800; op = 110;
#30 a = 29358; b = 22431; op = 110;
#30 a = 27440; b = 23793; op = 110;
#30 a = 7240; b = 38611; op = 110;
#30 a = 56; b = 13804; op = 110;
#30 a = 18273; b = 1061; op = 110;
#30 a = 54842; b = 19418; op = 110;
#30 a = 56626; b = 51259; op = 110;
#30 a = 27550; b = 8497; op = 110;
#30 a = 5238; b = 12278; op = 110;
#30 a = 49221; b = 56535; op = 110;
#30 a = 59290; b = 10715; op = 110;
#30 a = 36359; b = 53204; op = 110;
#30 a = 368; b = 12734; op = 110;
#30 a = 11957; b = 53170; op = 110;
#30 a = 37603; b = 34573; op = 110;
#30 a = 52925; b = 45044; op = 110;
#30 a = 20709; b = 41270; op = 110;
#30 a = 18155; b = 1680; op = 110;
#30 a = 18660; b = 4086; op = 110;
#30 a = 11276; b = 43946; op = 110;
#30 a = 18332; b = 31551; op = 110;
#30 a = 29710; b = 20079; op = 110;
#30 a = 35270; b = 48229; op = 110;
#30 a = 53156; b = 18795; op = 110;
#30 a = 54093; b = 44742; op = 110;
#30 a = 27206; b = 36711; op = 110;
#30 a = 4865; b = 8372; op = 110;
#30 a = 48405; b = 23458; op = 110;
#30 a = 44100; b = 54624; op = 110;
#30 a = 42107; b = 58571; op = 110;
#30 a = 12802; b = 18148; op = 110;
#30 a = 33809; b = 11864; op = 110;
#30 a = 22367; b = 49612; op = 110;
#30 a = 7258; b = 26182; op = 110;
#30 a = 32360; b = 56290; op = 110;
#30 a = 15149; b = 36590; op = 110;
#30 a = 40779; b = 24246; op = 110;
#30 a = 47952; b = 19872; op = 110;
#30 a = 37602; b = 4006; op = 110;
#30 a = 47583; b = 31711; op = 110;
#30 a = 39658; b = 49807; op = 110;
#30 a = 31468; b = 7545; op = 110;
#30 a = 58546; b = 36144; op = 110;
#30 a = 59233; b = 33793; op = 110;
#30 a = 54031; b = 44920; op = 110;
#30 a = 15649; b = 1162; op = 110;
#30 a = 47628; b = 19308; op = 110;
#30 a = 39564; b = 37794; op = 110;
#30 a = 36159; b = 1910; op = 110;
#30 a = 51617; b = 14632; op = 110;
#30 a = 59223; b = 42220; op = 110;
#30 a = 14909; b = 43052; op = 110;
#30 a = 20401; b = 24508; op = 110;
#30 a = 32962; b = 41154; op = 110;
#30 a = 48554; b = 8466; op = 110;
#30 a = 27732; b = 1571; op = 110;
#30 a = 15567; b = 21254; op = 110;
#30 a = 1180; b = 15040; op = 110;
#30 a = 26960; b = 53765; op = 110;
#30 a = 56399; b = 25475; op = 110;
#30 a = 36691; b = 20666; op = 110;
#30 a = 53929; b = 20676; op = 110;
#30 a = 21700; b = 34296; op = 110;
#30 a = 4435; b = 25892; op = 110;
#30 a = 2826; b = 20167; op = 110;
#30 a = 12644; b = 28650; op = 110;
#30 a = 20501; b = 49288; op = 110;
#30 a = 14947; b = 17848; op = 110;
#30 a = 43411; b = 56935; op = 110;
#30 a = 36586; b = 19945; op = 110;
#30 a = 33763; b = 52764; op = 110;
#30 a = 41606; b = 20105; op = 110;
#30 a = 54817; b = 12286; op = 110;
#30 a = 58299; b = 3345; op = 110;
#30 a = 607; b = 12357; op = 110;
#30 a = 11813; b = 3325; op = 110;
#30 a = 28404; b = 44314; op = 110;
#30 a = 21881; b = 58700; op = 110;
#30 a = 19054; b = 31965; op = 110;
#30 a = 56553; b = 40628; op = 110;
#30 a = 56900; b = 4722; op = 110;
#30 a = 29287; b = 33471; op = 110;
#30 a = 2406; b = 41098; op = 110;
#30 a = 48929; b = 58661; op = 110;
#30 a = 1686; b = 52745; op = 110;
#30 a = 3850; b = 50952; op = 110;
#30 a = 56143; b = 53881; op = 110;
#30 a = 57274; b = 29734; op = 110;
#30 a = 4931; b = 27339; op = 110;
#30 a = 11243; b = 4191; op = 110;
#30 a = 30404; b = 39269; op = 110;
#30 a = 31236; b = 4739; op = 110;
#30 a = 24024; b = 33548; op = 110;
#30 a = 17587; b = 22326; op = 110;
#30 a = 46159; b = 16079; op = 110;
#30 a = 38771; b = 58596; op = 110;
#30 a = 39504; b = 42733; op = 110;
#30 a = 35022; b = 40187; op = 110;
#30 a = 879; b = 28613; op = 110;
#30 a = 58971; b = 48873; op = 110;
#30 a = 11323; b = 2968; op = 110;
#30 a = 26344; b = 14419; op = 110;
#30 a = 47157; b = 20893; op = 110;
#30 a = 11027; b = 16430; op = 110;
#30 a = 39259; b = 15329; op = 110;
#30 a = 6194; b = 56382; op = 110;
#30 a = 8833; b = 45560; op = 110;
#30 a = 11154; b = 10985; op = 110;
#30 a = 29825; b = 49573; op = 110;
#30 a = 37629; b = 49719; op = 110;
#30 a = 17418; b = 32833; op = 110;
#30 a = 24885; b = 15401; op = 110;
#30 a = 39956; b = 6860; op = 110;
#30 a = 11741; b = 28947; op = 110;
#30 a = 49299; b = 27597; op = 110;
#30 a = 22006; b = 16790; op = 110;
#30 a = 57225; b = 20999; op = 110;
#30 a = 46054; b = 1342; op = 110;
#30 a = 38358; b = 1019; op = 110;
#30 a = 18070; b = 47765; op = 110;
#30 a = 42571; b = 9300; op = 110;
#30 a = 24306; b = 37283; op = 110;
#30 a = 39677; b = 14195; op = 110;
#30 a = 39155; b = 31779; op = 110;
#30 a = 756; b = 27575; op = 110;
#30 a = 52985; b = 30371; op = 110;
#30 a = 39043; b = 56360; op = 110;
#30 a = 11314; b = 42967; op = 110;
#30 a = 49874; b = 13409; op = 110;
#30 a = 34808; b = 5882; op = 110;
#30 a = 52726; b = 18488; op = 110;
#30 a = 19638; b = 42850; op = 110;
#30 a = 51171; b = 45419; op = 110;
#30 a = 25962; b = 36862; op = 110;
#30 a = 13048; b = 21992; op = 110;
#30 a = 58758; b = 1359; op = 110;
#30 a = 9144; b = 53048; op = 110;
#30 a = 19377; b = 18817; op = 110;
#30 a = 30457; b = 23594; op = 110;
#30 a = 27083; b = 55909; op = 110;
#30 a = 43733; b = 25656; op = 110;
#30 a = 15309; b = 47148; op = 110;
#30 a = 13118; b = 28760; op = 110;
#30 a = 27822; b = 22882; op = 110;
#30 a = 57039; b = 30817; op = 110;
#30 a = 44195; b = 8292; op = 110;
#30 a = 28733; b = 25368; op = 110;
#30 a = 44510; b = 16351; op = 110;
#30 a = 17676; b = 46902; op = 110;
#30 a = 16503; b = 29191; op = 110;
#30 a = 38206; b = 43255; op = 110;
#30 a = 40200; b = 49456; op = 110;
#30 a = 33254; b = 21442; op = 110;
#30 a = 19537; b = 6413; op = 110;
#30 a = 49819; b = 51888; op = 110;
#30 a = 15004; b = 20547; op = 110;
#30 a = 59880; b = 12283; op = 110;
#30 a = 2684; b = 25736; op = 110;
#30 a = 43680; b = 41764; op = 110;
#30 a = 1806; b = 12062; op = 110;
#30 a = 9870; b = 51105; op = 110;
#30 a = 19490; b = 27206; op = 110;
#30 a = 16651; b = 50209; op = 110;
#30 a = 37459; b = 47330; op = 110;
#30 a = 20649; b = 22558; op = 110;
#30 a = 50672; b = 29676; op = 110;
#30 a = 14764; b = 34430; op = 110;
#30 a = 20575; b = 4844; op = 110;
#30 a = 50392; b = 12997; op = 110;
#30 a = 31160; b = 11514; op = 110;
#30 a = 2214; b = 54778; op = 110;
#30 a = 44301; b = 57424; op = 110;
#30 a = 14576; b = 41268; op = 110;
#30 a = 17641; b = 58827; op = 110;
#30 a = 41227; b = 7265; op = 110;
#30 a = 12694; b = 42686; op = 110;
#30 a = 28949; b = 48020; op = 110;
#30 a = 26393; b = 58195; op = 110;
#30 a = 13284; b = 49609; op = 110;
#30 a = 26456; b = 42559; op = 110;
#30 a = 59710; b = 39765; op = 110;
#30 a = 5947; b = 29089; op = 110;
#30 a = 58983; b = 26255; op = 110;
#30 a = 1648; b = 24663; op = 110;
#30 a = 34548; b = 40052; op = 110;
#30 a = 57865; b = 10684; op = 110;
#30 a = 45630; b = 5852; op = 110;
#30 a = 52512; b = 46882; op = 110;
#30 a = 31858; b = 23511; op = 110;
#30 a = 30202; b = 4744; op = 110;
#30 a = 70; b = 16899; op = 110;
#30 a = 52489; b = 41624; op = 110;
#30 a = 45510; b = 12878; op = 110;
#30 a = 3564; b = 33216; op = 110;
#30 a = 42572; b = 36098; op = 110;
#30 a = 49169; b = 43978; op = 110;
#30 a = 12590; b = 27569; op = 110;
#30 a = 20123; b = 26938; op = 110;
#30 a = 44049; b = 15966; op = 110;
#30 a = 20222; b = 53796; op = 110;
#30 a = 44316; b = 45542; op = 110;
#30 a = 47015; b = 31112; op = 110;
#30 a = 46759; b = 30505; op = 110;
#30 a = 48121; b = 59723; op = 110;
#30 a = 20402; b = 55321; op = 110;
#30 a = 58578; b = 35411; op = 110;
#30 a = 25042; b = 56030; op = 110;
#30 a = 7372; b = 35071; op = 110;
#30 a = 8870; b = 47779; op = 110;
#30 a = 2591; b = 15168; op = 110;
#30 a = 776; b = 9120; op = 110;
#30 a = 20964; b = 20311; op = 110;
#30 a = 32863; b = 28389; op = 110;
#30 a = 52340; b = 29837; op = 110;
#30 a = 12784; b = 45280; op = 110;
#30 a = 7918; b = 27913; op = 110;
#30 a = 14261; b = 42892; op = 110;
#30 a = 31448; b = 9745; op = 110;
#30 a = 48134; b = 9622; op = 110;
#30 a = 38173; b = 50465; op = 110;
#30 a = 16436; b = 30796; op = 110;
#30 a = 42069; b = 641; op = 110;
#30 a = 32949; b = 41125; op = 110;
#30 a = 56386; b = 25510; op = 110;
#30 a = 26233; b = 5703; op = 110;
#30 a = 6678; b = 17255; op = 110;
#30 a = 53851; b = 10585; op = 110;
#30 a = 10162; b = 26522; op = 110;
#30 a = 39027; b = 4581; op = 110;
#30 a = 10730; b = 53579; op = 110;
#30 a = 52328; b = 25513; op = 110;
#30 a = 22596; b = 14328; op = 110;
#30 a = 7811; b = 18875; op = 110;
#30 a = 56799; b = 844; op = 110;
#30 a = 45534; b = 45911; op = 110;
#30 a = 1104; b = 40278; op = 110;
#30 a = 20123; b = 16198; op = 110;
#30 a = 35399; b = 43525; op = 110;
#30 a = 59602; b = 48012; op = 110;
#30 a = 43888; b = 40930; op = 110;
#30 a = 42242; b = 814; op = 110;
#30 a = 49621; b = 41290; op = 110;
#30 a = 32105; b = 42911; op = 110;
#30 a = 29569; b = 16583; op = 110;
#30 a = 15407; b = 8966; op = 110;
#30 a = 37824; b = 23594; op = 110;
#30 a = 30876; b = 49773; op = 110;
#30 a = 35267; b = 34279; op = 110;
#30 a = 38921; b = 8647; op = 110;
#30 a = 4063; b = 812; op = 110;
#30 a = 8308; b = 12831; op = 110;
#30 a = 54293; b = 5919; op = 110;
#30 a = 30765; b = 39322; op = 110;
#30 a = 40652; b = 17684; op = 110;
#30 a = 58061; b = 21769; op = 110;
#30 a = 23673; b = 5672; op = 110;
#30 a = 58343; b = 27277; op = 110;
#30 a = 8097; b = 26333; op = 110;
#30 a = 38807; b = 9638; op = 110;
#30 a = 53493; b = 49489; op = 110;
#30 a = 29814; b = 42906; op = 110;
#30 a = 13660; b = 17213; op = 110;
#30 a = 30992; b = 6879; op = 110;
#30 a = 59727; b = 37608; op = 110;
#30 a = 49996; b = 2917; op = 110;
#30 a = 46942; b = 43078; op = 110;
#30 a = 55242; b = 55107; op = 110;
#30 a = 39664; b = 34576; op = 110;
#30 a = 24396; b = 39100; op = 110;
#30 a = 29703; b = 51841; op = 110;
#30 a = 51531; b = 30061; op = 110;
#30 a = 56738; b = 36234; op = 110;
#30 a = 48234; b = 50167; op = 110;
#30 a = 32348; b = 27218; op = 110;
#30 a = 25383; b = 5955; op = 110;
#30 a = 52914; b = 21166; op = 110;
#30 a = 55726; b = 49303; op = 110;
#30 a = 58401; b = 24185; op = 110;
#30 a = 23080; b = 4243; op = 110;
#30 a = 21197; b = 2512; op = 110;
#30 a = 25744; b = 5416; op = 110;
#30 a = 49695; b = 24973; op = 110;
#30 a = 39014; b = 35606; op = 110;
#30 a = 18342; b = 48477; op = 110;
#30 a = 17629; b = 50080; op = 110;
#30 a = 33438; b = 58144; op = 110;
#30 a = 17455; b = 54607; op = 110;
#30 a = 48142; b = 36701; op = 110;
#30 a = 22064; b = 30431; op = 110;
#30 a = 35723; b = 55999; op = 110;
#30 a = 23967; b = 42730; op = 110;
#30 a = 32378; b = 22576; op = 110;
#30 a = 13113; b = 14895; op = 110;
#30 a = 12659; b = 43729; op = 110;
#30 a = 8136; b = 59647; op = 110;
#30 a = 4033; b = 34867; op = 110;
#30 a = 46937; b = 31556; op = 110;
#30 a = 38150; b = 33717; op = 110;
#30 a = 57003; b = 8270; op = 110;
#30 a = 10779; b = 24474; op = 110;
#30 a = 52003; b = 5371; op = 110;
#30 a = 6740; b = 36998; op = 110;
#30 a = 55325; b = 49729; op = 110;
#30 a = 51970; b = 48437; op = 110;
#30 a = 21437; b = 3707; op = 110;
#30 a = 49907; b = 40696; op = 110;
#30 a = 52067; b = 29391; op = 110;
#30 a = 34228; b = 47245; op = 110;
#30 a = 956; b = 36664; op = 110;
#30 a = 13686; b = 12537; op = 110;
#30 a = 31733; b = 1973; op = 110;
#30 a = 54926; b = 36389; op = 110;
#30 a = 58347; b = 50221; op = 110;
#30 a = 11095; b = 47923; op = 110;
#30 a = 1502; b = 44701; op = 110;
#30 a = 45938; b = 50555; op = 110;
#30 a = 26340; b = 49055; op = 110;
#30 a = 42285; b = 14566; op = 110;
#30 a = 20281; b = 22552; op = 110;
#30 a = 15394; b = 21158; op = 110;
#30 a = 1268; b = 11295; op = 110;
#30 a = 16982; b = 59664; op = 110;
#30 a = 36469; b = 26789; op = 110;
#30 a = 48194; b = 3095; op = 110;
#30 a = 24891; b = 44709; op = 110;
#30 a = 25614; b = 49190; op = 110;
#30 a = 37970; b = 28266; op = 110;
#30 a = 6937; b = 10490; op = 110;
#30 a = 12809; b = 13911; op = 110;
#30 a = 19413; b = 218; op = 110;
#30 a = 18306; b = 28695; op = 110;
#30 a = 46768; b = 32052; op = 110;
#30 a = 31618; b = 23426; op = 110;
#30 a = 38221; b = 29621; op = 110;
#30 a = 51368; b = 5832; op = 110;
#30 a = 25425; b = 52740; op = 110;
#30 a = 38811; b = 10525; op = 110;
#30 a = 54745; b = 35035; op = 110;
#30 a = 47387; b = 2561; op = 110;
#30 a = 22792; b = 28419; op = 110;
#30 a = 14650; b = 27467; op = 110;
#30 a = 54751; b = 58700; op = 110;
#30 a = 34788; b = 47729; op = 110;
#30 a = 2533; b = 9670; op = 110;
#30 a = 35128; b = 10263; op = 110;
#30 a = 29254; b = 47966; op = 110;
#30 a = 20923; b = 46065; op = 110;
#30 a = 22968; b = 7352; op = 110;
#30 a = 37250; b = 32855; op = 110;
#30 a = 54520; b = 53062; op = 110;
#30 a = 41805; b = 16068; op = 110;
#30 a = 20179; b = 46882; op = 110;
#30 a = 7764; b = 20938; op = 110;
#30 a = 44129; b = 14478; op = 110;
#30 a = 22777; b = 38231; op = 110;
#30 a = 20331; b = 12037; op = 110;
#30 a = 43932; b = 7996; op = 110;
#30 a = 55149; b = 24413; op = 110;
#30 a = 1133; b = 51231; op = 110;
#30 a = 12183; b = 58844; op = 110;
#30 a = 20092; b = 45567; op = 110;
#30 a = 29293; b = 52404; op = 110;
#30 a = 29517; b = 4415; op = 110;
#30 a = 14639; b = 2493; op = 110;
#30 a = 50952; b = 22610; op = 110;
#30 a = 32531; b = 7597; op = 110;
#30 a = 47692; b = 24257; op = 110;
#30 a = 15533; b = 23030; op = 110;
#30 a = 1315; b = 22555; op = 110;
#30 a = 49872; b = 28508; op = 110;
#30 a = 44657; b = 2458; op = 110;
#30 a = 4655; b = 53937; op = 110;
#30 a = 25478; b = 47886; op = 110;
#30 a = 12060; b = 21807; op = 110;
#30 a = 28883; b = 45992; op = 110;
#30 a = 53714; b = 21970; op = 110;
#30 a = 39513; b = 58725; op = 110;
#30 a = 31086; b = 20464; op = 110;
#30 a = 31005; b = 17269; op = 110;
#30 a = 34040; b = 27957; op = 110;
#30 a = 15415; b = 39719; op = 110;
#30 a = 15776; b = 16575; op = 110;
#30 a = 24138; b = 57331; op = 110;
#30 a = 56419; b = 46034; op = 110;
#30 a = 16622; b = 31715; op = 110;
#30 a = 25196; b = 57881; op = 110;
#30 a = 20201; b = 25087; op = 110;
#30 a = 52375; b = 42939; op = 110;
#30 a = 14108; b = 18835; op = 110;
#30 a = 41073; b = 55990; op = 110;
#30 a = 30521; b = 24703; op = 110;
#30 a = 56283; b = 6490; op = 110;
#30 a = 14323; b = 23548; op = 110;
#30 a = 35405; b = 44068; op = 110;
#30 a = 27534; b = 34374; op = 110;
#30 a = 45528; b = 23413; op = 110;
#30 a = 341; b = 1482; op = 110;
#30 a = 57604; b = 34735; op = 110;
#30 a = 32522; b = 1293; op = 110;
#30 a = 16088; b = 2668; op = 110;
#30 a = 15512; b = 58198; op = 110;
#30 a = 51479; b = 58298; op = 110;
#30 a = 45764; b = 24761; op = 110;
#30 a = 24263; b = 9303; op = 110;
#30 a = 46722; b = 43489; op = 110;
#30 a = 52430; b = 15685; op = 110;
#30 a = 57796; b = 21849; op = 110;
#30 a = 5109; b = 5546; op = 110;
#30 a = 6509; b = 28792; op = 110;
#30 a = 718; b = 36710; op = 110;
#30 a = 5988; b = 16487; op = 110;
#30 a = 38194; b = 51954; op = 110;
#30 a = 5988; b = 49679; op = 110;
#30 a = 39267; b = 31762; op = 110;
#30 a = 26128; b = 9764; op = 110;
#30 a = 7312; b = 45046; op = 110;
#30 a = 35812; b = 1672; op = 110;
#30 a = 3831; b = 20723; op = 110;
#30 a = 10150; b = 18973; op = 110;
#30 a = 21892; b = 50713; op = 110;
#30 a = 50267; b = 42187; op = 110;
#30 a = 43736; b = 3632; op = 110;
#30 a = 42487; b = 4330; op = 110;
#30 a = 5413; b = 16244; op = 110;
#30 a = 37996; b = 24781; op = 110;
#30 a = 55766; b = 38314; op = 110;
#30 a = 8707; b = 3627; op = 110;
#30 a = 3979; b = 9566; op = 110;
#30 a = 45481; b = 50667; op = 110;
#30 a = 18369; b = 50459; op = 110;
#30 a = 23264; b = 55851; op = 110;
#30 a = 48976; b = 4549; op = 110;
#30 a = 24183; b = 40365; op = 110;
#30 a = 17071; b = 18071; op = 110;
#30 a = 11764; b = 24159; op = 110;
#30 a = 55250; b = 58740; op = 110;
#30 a = 4909; b = 32613; op = 110;
#30 a = 54195; b = 39820; op = 110;
#30 a = 24630; b = 41990; op = 110;
#30 a = 39823; b = 19341; op = 110;
#30 a = 14772; b = 7631; op = 110;
#30 a = 38055; b = 13859; op = 110;
#30 a = 28880; b = 11335; op = 110;
#30 a = 37414; b = 40462; op = 110;
#30 a = 648; b = 8337; op = 110;
#30 a = 29634; b = 37726; op = 110;
#30 a = 27807; b = 40375; op = 110;
#30 a = 49884; b = 45486; op = 110;
#30 a = 16052; b = 24474; op = 110;
#30 a = 32066; b = 47514; op = 110;
#30 a = 49585; b = 56339; op = 110;
#30 a = 23028; b = 53150; op = 110;
#30 a = 45978; b = 28068; op = 110;
#30 a = 36419; b = 8428; op = 110;
#30 a = 11781; b = 8928; op = 110;
#30 a = 4981; b = 5801; op = 110;
#30 a = 39849; b = 59251; op = 110;
#30 a = 10918; b = 56517; op = 110;
#30 a = 45262; b = 22287; op = 110;
#30 a = 35560; b = 36694; op = 110;
#30 a = 23780; b = 17557; op = 110;
#30 a = 45099; b = 2992; op = 110;
#30 a = 22768; b = 47196; op = 110;
#30 a = 7959; b = 3715; op = 110;
#30 a = 49761; b = 20033; op = 110;
#30 a = 17206; b = 50096; op = 110;
#30 a = 26145; b = 56396; op = 110;
#30 a = 21999; b = 38569; op = 110;
#30 a = 3015; b = 26874; op = 110;
#30 a = 5997; b = 33957; op = 110;
#30 a = 34921; b = 22828; op = 110;
#30 a = 17982; b = 17596; op = 110;
#30 a = 18638; b = 8588; op = 110;
#30 a = 35543; b = 55621; op = 110;
#30 a = 48865; b = 56855; op = 110;
#30 a = 35925; b = 10922; op = 110;
#30 a = 51170; b = 23307; op = 110;
#30 a = 21214; b = 14724; op = 110;
#30 a = 38455; b = 20174; op = 110;
#30 a = 41382; b = 50425; op = 110;
#30 a = 31456; b = 26584; op = 110;
#30 a = 4686; b = 16782; op = 110;
#30 a = 55272; b = 23199; op = 110;
#30 a = 21766; b = 39818; op = 110;
#30 a = 53943; b = 58525; op = 110;
#30 a = 45107; b = 44714; op = 110;
#30 a = 26341; b = 31424; op = 110;
#30 a = 18348; b = 8090; op = 110;
#30 a = 22344; b = 32173; op = 110;
#30 a = 30750; b = 12662; op = 110;
#30 a = 27214; b = 6194; op = 110;
#30 a = 3504; b = 20765; op = 110;
#30 a = 31622; b = 14631; op = 110;
#30 a = 58080; b = 40879; op = 110;
#30 a = 39193; b = 52768; op = 110;
#30 a = 14988; b = 995; op = 110;
#30 a = 32310; b = 30706; op = 110;
#30 a = 49101; b = 28296; op = 110;
#30 a = 27243; b = 38527; op = 110;
#30 a = 12254; b = 28790; op = 110;
#30 a = 49040; b = 57312; op = 110;
#30 a = 11066; b = 5487; op = 110;
#30 a = 3229; b = 16974; op = 110;
#30 a = 21731; b = 5719; op = 110;
#30 a = 40123; b = 19692; op = 110;
#30 a = 42207; b = 49421; op = 110;
#30 a = 38680; b = 57109; op = 110;
#30 a = 10525; b = 53605; op = 110;
#30 a = 23092; b = 8061; op = 110;
#30 a = 47350; b = 23780; op = 110;
#30 a = 4633; b = 51975; op = 110;
#30 a = 45774; b = 36183; op = 110;
#30 a = 5671; b = 44419; op = 110;
#30 a = 6521; b = 59504; op = 110;
#30 a = 15181; b = 16321; op = 110;
#30 a = 54810; b = 19039; op = 110;
#30 a = 8276; b = 18231; op = 110;
#30 a = 42695; b = 12041; op = 110;
#30 a = 14997; b = 42474; op = 110;
#30 a = 54568; b = 13607; op = 110;
#30 a = 23723; b = 58844; op = 110;
#30 a = 10335; b = 18717; op = 110;
#30 a = 53443; b = 28499; op = 110;
#30 a = 34369; b = 8245; op = 110;
#30 a = 42544; b = 20450; op = 110;
#30 a = 5090; b = 27991; op = 110;
#30 a = 443; b = 49494; op = 110;
#30 a = 7567; b = 19336; op = 110;
#30 a = 45591; b = 30143; op = 110;
#30 a = 10197; b = 41245; op = 110;
#30 a = 26034; b = 29145; op = 110;
#30 a = 27807; b = 40986; op = 110;
#30 a = 11976; b = 29430; op = 110;
#30 a = 44188; b = 5867; op = 110;
#30 a = 23602; b = 15882; op = 110;
#30 a = 34911; b = 30717; op = 110;
#30 a = 37372; b = 15922; op = 110;
#30 a = 31296; b = 47162; op = 110;
#30 a = 11955; b = 8641; op = 110;
#30 a = 42656; b = 928; op = 110;
#30 a = 38397; b = 27497; op = 110;
#30 a = 15082; b = 57213; op = 110;
#30 a = 20067; b = 56290; op = 110;
#30 a = 52788; b = 9577; op = 110;
#30 a = 17993; b = 57947; op = 110;
#30 a = 6885; b = 33984; op = 110;
#30 a = 41855; b = 48026; op = 110;
#30 a = 8560; b = 43067; op = 110;
#30 a = 1328; b = 35985; op = 110;
#30 a = 12351; b = 50633; op = 110;
#30 a = 439; b = 30527; op = 110;
#30 a = 1643; b = 25295; op = 110;
#30 a = 54609; b = 10528; op = 110;
#30 a = 9383; b = 13497; op = 110;
#30 a = 13549; b = 11347; op = 110;
#30 a = 18397; b = 6204; op = 110;
#30 a = 32672; b = 55334; op = 110;
#30 a = 42480; b = 5930; op = 110;
#30 a = 21270; b = 49791; op = 110;
#30 a = 13377; b = 31024; op = 110;
#30 a = 20515; b = 2057; op = 110;
#30 a = 24396; b = 24335; op = 110;
#30 a = 36727; b = 17753; op = 110;
#30 a = 47986; b = 46197; op = 110;
#30 a = 4911; b = 20221; op = 110;
#30 a = 59570; b = 12536; op = 110;
#30 a = 7048; b = 25440; op = 110;
#30 a = 15281; b = 7951; op = 110;
#30 a = 53071; b = 51292; op = 110;
#30 a = 42489; b = 2317; op = 110;
#30 a = 4308; b = 43900; op = 110;
#30 a = 32317; b = 36731; op = 110;
#30 a = 54653; b = 23469; op = 110;
#30 a = 14394; b = 34672; op = 110;
#30 a = 10103; b = 30017; op = 110;
#30 a = 55288; b = 56079; op = 110;
#30 a = 47687; b = 58719; op = 110;
#30 a = 34096; b = 24350; op = 110;
#30 a = 49278; b = 30954; op = 110;
#30 a = 5225; b = 7838; op = 110;
#30 a = 491; b = 42540; op = 110;
#30 a = 1787; b = 40588; op = 110;
#30 a = 1450; b = 34559; op = 110;
#30 a = 50676; b = 17171; op = 110;
#30 a = 16346; b = 38425; op = 110;
#30 a = 234; b = 19; op = 110;
$display($time,, "a=%d, b=%d, s=%d, cout=%b, op=%b, choice=%b, q=%d", a, b, s, cout, op, choice, q);
end
endmodule
